/**
 * $Id: red_pitaya_top.v 1271 2014-02-25 12:32:34Z matej.oblak $
 *
 * @brief Red Pitaya TOP module. It connects external pins and PS part with 
 *        other application modules. 
 *
 * @Author Matej Oblak
 *
 * (c) Red Pitaya  http://www.redpitaya.com
 *
 * This part of code is written in Verilog hardware description language (HDL).
 * Please visit http://en.wikipedia.org/wiki/Verilog
 * for more details on the language used herein.
 */


/**
 * GENERAL DESCRIPTION:
 *
 * Top module connects PS part with rest of Red Pitaya applications.  
 *
 *
 *                   /-------\      
 *   PS DDR <------> |  PS   |      AXI <-> custom bus
 *   PS MIO <------> |   /   | <------------+
 *   PS CLK -------> |  ARM  |              |
 *                   \-------/              |
 *                                          |
 *                            /-------\     |
 *                         -> | SCOPE | <---+
 *                         |  \-------/     |
 *                         |                |
 *            /--------\   |   /-----\      |
 *   ADC ---> |        | --+-> |     |      |
 *            | ANALOG |       | PID | <----+
 *   DAC <--- |        | <---- |     |      |
 *            \--------/   ^   \-----/      |
 *                         |                |
 *                         |  /-------\     |
 *                         -- |  ASG  | <---+ 
 *                            \-------/     |
 *                                          |
 *             /--------\                   |
 *    RX ----> |        |                   |
 *   SATA      | DAISY  | <-----------------+
 *    TX <---- |        | 
 *             \--------/ 
 *               |    |
 *               |    |
 *               (FREE)
 *
 *
 * Inside the analog module, ADC data is translated from unsigned neg-slope into
 * two's complement. Similar is done on DAC data.
 *
 * Scope module stores data from ADC into RAM, arbitrary signal generator (ASG)
 * sends data from RAM to DAC. MIMO PID uses ADC ADC as input and DAC as its output.
 *
 * Daisy chain connects with other boards with fast serial link. Data which is
 * sent and received is at the moment undefined. This is left for the user.
 * 
 */

module red_pitaya_top (
   // PS connections
   inout  [54-1: 0] FIXED_IO_mio       ,
   inout            FIXED_IO_ps_clk    ,
   inout            FIXED_IO_ps_porb   ,
   inout            FIXED_IO_ps_srstb  ,
   inout            FIXED_IO_ddr_vrn   ,
   inout            FIXED_IO_ddr_vrp   ,
   // DDR
   inout  [15-1: 0] DDR_addr           ,
   inout  [ 3-1: 0] DDR_ba             ,
   inout            DDR_cas_n          ,
   inout            DDR_ck_n           ,
   inout            DDR_ck_p           ,
   inout            DDR_cke            ,
   inout            DDR_cs_n           ,
   inout  [ 4-1: 0] DDR_dm             ,
   inout  [32-1: 0] DDR_dq             ,
   inout  [ 4-1: 0] DDR_dqs_n          ,
   inout  [ 4-1: 0] DDR_dqs_p          ,
   inout            DDR_odt            ,
   inout            DDR_ras_n          ,
   inout            DDR_reset_n        ,
   inout            DDR_we_n           ,

   // Red Pitaya periphery
  
   // ADC
   input  [16-1: 2] adc_dat_a_i        ,  // ADC CH1
   input  [16-1: 2] adc_dat_b_i        ,  // ADC CH2
   input            adc_clk_p_i        ,  // ADC data clock
   input            adc_clk_n_i        ,  // ADC data clock
   output [ 2-1: 0] adc_clk_o          ,  // optional ADC clock source
   output           adc_cdcs_o         ,  // ADC clock duty cycle stabilizer
   // DAC
   output [14-1: 0] dac_dat_o          ,  // DAC combined data
   output           dac_wrt_o          ,  // DAC write
   output           dac_sel_o          ,  // DAC channel select
   output           dac_clk_o          ,  // DAC clock
   output           dac_rst_o          ,  // DAC reset
   // PWM DAC
   output [ 4-1: 0] dac_pwm_o          ,  // serial PWM DAC
   // XADC
   input  [ 5-1: 0] vinp_i             ,  // voltages p
   input  [ 5-1: 0] vinn_i             ,  // voltages n
   // Expansion connector
   inout  [ 8-1: 0] exp_p_io           ,
   inout  [ 8-1: 0] exp_n_io           ,
   // SATA connector
   output [ 2-1: 0] daisy_p_o          ,  // line 1 is clock capable
   output [ 2-1: 0] daisy_n_o          ,
   input  [ 2-1: 0] daisy_p_i          ,  // line 1 is clock capable
   input  [ 2-1: 0] daisy_n_i          ,
   // LED
   output [ 8-1: 0] led_o       
);


localparam       SMC = 8                     ;  // Sub Module Count

//---------------------------------------------------------------------------------
//
//  Connections to PS

wire  [  4-1: 0] fclk                        ;  //[0] = 125 MHz, [1] = 250 MHz, [2] = 50 MHz, [3] = 200 MHz  based on PS connected oscillator
wire  [  4-1: 0] frstn                       ;

wire             ps_sys_clk                  ;
wire             ps_sys_rstn                 ;
wire  [ 32-1: 0] ps_sys_addr                 ;
wire  [ 32-1: 0] ps_sys_wdata                ;
wire  [  4-1: 0] ps_sys_sel                  ;
wire             ps_sys_wen                  ;
wire             ps_sys_ren                  ;
wire  [ 32-1: 0] ps_sys_rdata                ;
wire             ps_sys_err                  ;
wire             ps_sys_ack                  ;

// AXI masters
wire             axi_clk    [1:0]            ;
wire             axi_rstn   [1:0]            ;
wire  [ 32-1: 0] axi_waddr  [1:0]            ;
wire  [ 64-1: 0] axi_wdata  [1:0]            ;
wire  [  8-1: 0] axi_wsel   [1:0]            ;
wire             axi_wvalid [1:0]            ;
wire  [  4-1: 0] axi_wlen   [1:0]            ;
wire             axi_wfixed [1:0]            ;
wire             axi_werr   [1:0]            ;
wire             axi_wrdy   [1:0]            ;


red_pitaya_ps i_ps (
  .FIXED_IO_mio     (FIXED_IO_mio     ),
  .FIXED_IO_ps_clk  (FIXED_IO_ps_clk  ),
  .FIXED_IO_ps_porb (FIXED_IO_ps_porb ),
  .FIXED_IO_ps_srstb(FIXED_IO_ps_srstb),
  .FIXED_IO_ddr_vrn (FIXED_IO_ddr_vrn ),
  .FIXED_IO_ddr_vrp (FIXED_IO_ddr_vrp ),
  // DDR
  .DDR_addr      (DDR_addr    ),
  .DDR_ba        (DDR_ba      ),
  .DDR_cas_n     (DDR_cas_n   ),
  .DDR_ck_n      (DDR_ck_n    ),
  .DDR_ck_p      (DDR_ck_p    ),
  .DDR_cke       (DDR_cke     ),
  .DDR_cs_n      (DDR_cs_n    ),
  .DDR_dm        (DDR_dm      ),
  .DDR_dq        (DDR_dq      ),
  .DDR_dqs_n     (DDR_dqs_n   ),
  .DDR_dqs_p     (DDR_dqs_p   ),
  .DDR_odt       (DDR_odt     ),
  .DDR_ras_n     (DDR_ras_n   ),
  .DDR_reset_n   (DDR_reset_n ),
  .DDR_we_n      (DDR_we_n    ),

  .fclk_clk_o    (fclk        ),
  .fclk_rstn_o   (frstn       ),
  // ADC analog inputs
  .vinp_i        (vinp_i      ),  // voltages p
  .vinn_i        (vinn_i      ),  // voltages n
   // system read/write channel
  .sys_clk_o     (ps_sys_clk  ),  // system clock
  .sys_rstn_o    (ps_sys_rstn ),  // system reset - active low
  .sys_addr_o    (ps_sys_addr ),  // system read/write address
  .sys_wdata_o   (ps_sys_wdata),  // system write data
  .sys_sel_o     (ps_sys_sel  ),  // system write byte select
  .sys_wen_o     (ps_sys_wen  ),  // system write enable
  .sys_ren_o     (ps_sys_ren  ),  // system read enable
  .sys_rdata_i   (ps_sys_rdata),  // system read data
  .sys_err_i     (ps_sys_err  ),  // system error indicator
  .sys_ack_i     (ps_sys_ack  ),  // system acknowledge signal
  // two AXI masters - concatenated
  .axi_clk_i     ( {axi_clk   [1], axi_clk   [0]} ),  // global clock
  .axi_rstn_i    ( {axi_rstn  [1], axi_rstn  [0]} ),  // global reset
  .axi_waddr_i   ( {axi_waddr [1], axi_waddr [0]} ),  // system write address
  .axi_wdata_i   ( {axi_wdata [1], axi_wdata [0]} ),  // system write data
  .axi_wsel_i    ( {axi_wsel  [1], axi_wsel  [0]} ),  // system write byte select
  .axi_wvalid_i  ( {axi_wvalid[1], axi_wvalid[0]} ),  // system write data valid
  .axi_wlen_i    ( {axi_wlen  [1], axi_wlen  [0]} ),  // system write burst length
  .axi_wfixed_i  ( {axi_wfixed[1], axi_wfixed[0]} ),  // system write burst type (fixed / incremental)
  .axi_werr_o    ( {axi_werr  [1], axi_werr  [0]} ),  // system write error
  .axi_wrdy_o    ( {axi_wrdy  [1], axi_wrdy  [0]} )    // system write ready
);

////////////////////////////////////////////////////////////////////////////////////////
// system bus decoder & multiplexer (it breaks memory addresses into SMC count regions)
////////////////////////////////////////////////////////////////////////////////////////

wire                sys_clk   = ps_sys_clk  ;
wire                sys_rstn  = ps_sys_rstn ;
wire  [    32-1: 0] sys_addr  = ps_sys_addr ;
wire  [    32-1: 0] sys_wdata = ps_sys_wdata;
wire  [     4-1: 0] sys_sel   = ps_sys_sel  ;
wire  [SMC   -1: 0] sys_wen                 ;
wire  [SMC   -1: 0] sys_ren                 ;
wire  [SMC*32-1: 0] sys_rdata               ;
wire  [SMC* 1-1: 0] sys_err                 ;
wire  [SMC* 1-1: 0] sys_ack                 ;
wire  [SMC   -1: 0] sys_cs                  ;

assign sys_cs = { {(SMC-1){1'b0}}, 1'h1 } << sys_addr[22:20] ;  // one-hot assignment

assign sys_wen = sys_cs & { SMC{ps_sys_wen} };
assign sys_ren = sys_cs & { SMC{ps_sys_ren} };

assign ps_sys_rdata = sys_rdata[sys_addr[22:20]*32+:32];

assign ps_sys_err   = |(sys_cs & sys_err);
assign ps_sys_ack   = |(sys_cs & sys_ack);


// unused system bus slave ports

assign sys_rdata[7*32+:32] = 32'h0; 
assign sys_err  [7       ] =  1'b0;
assign sys_ack  [7       ] =  1'b1;


////////////////////////////////////////////////////////////////////////////////
// local signals
////////////////////////////////////////////////////////////////////////////////

// PLL signals
wire                  clk_adc_125mhz_000deg;
wire                  clk_adc_250mhz_000deg;
wire                  clk_adc_250mhz_315deg;
wire                  clk_adc_200mhz_000deg;
wire                  clk_adc_20mhz_000deg;
wire                  pll_locked;

// PWM reset
reg                   pwm_rstn;

// ADC signals
reg                   adc_rstn;
reg          [14-1:0] adc_dat_a, adc_dat_b;
wire  signed [14-1:0] adc_a    , adc_b    ;

// DAC signals
//wire                dac_clk_1x;
//wire                dac_clk_2x;
//wire                dac_clk_2p;
reg                   dac_rst;
reg          [14-1:0] dac_dat_a, dac_dat_b;
wire         [14-1:0] dac_a    , dac_b    ;
wire  signed [15-1:0] dac_a_sum, dac_b_sum;

// ASG
wire  signed [14-1:0] asg_a    , asg_b    ;

// PID
wire  signed [14-1:0] pid_a    , pid_b    ;

// configuration
wire                  digital_loop;


////////////////////////////////////////////////////////////////////////////////
// PLL (clock and reset)
////////////////////////////////////////////////////////////////////////////////

clk_adc_pll i_clk_adc_pll (
  // Status and control signals
  .rstn                     ( frstn[0]              ),
  .pll_locked               ( pll_locked            ),

 // Clock in ports
  .adc_clk_i_p              ( adc_clk_p_i           ),
  .adc_clk_i_n              ( adc_clk_n_i           ),

  // Clock out ports
  .clk_adc_125mhz_000deg    ( clk_adc_125mhz_000deg ),
  .clk_adc_250mhz_000deg    ( clk_adc_250mhz_000deg ),
  .clk_adc_250mhz_315deg    ( clk_adc_250mhz_315deg ),
  .clk_adc_200mhz_000deg    ( clk_adc_200mhz_000deg ),
  .clk_adc_20mhz_000deg     ( clk_adc_20mhz_000deg  )
);

/*
// differential clock input
IBUFDS i_clk (.I (adc_clk_p_i), .IB (adc_clk_n_i), .O (adc_clk_in));  // differential clock input

red_pitaya_pll i_pll (
  // inputs
  .clk         (adc_clk_in),  // clock
  .rstn        (frstn[0]  ),  // reset - active low
  // output clocks
  .clk_adc     (pll_adc_clk   ),  // ADC clock
  .clk_dac_1x  (pll_dac_clk_1x),  // DAC clock 125MHz
  .clk_dac_2x  (pll_dac_clk_2x),  // DAC clock 250MHz
  .clk_dac_2p  (pll_dac_clk_2p),  // DAC clock 250MHz -45DGR
  .clk_ser     (pll_ser_clk   ),  // fast serial clock 200MHz
  .clk_pwm     (pll_pwm_clk   ),  // PWM clock
  // status outputs
  .pll_locked  (pll_locked)
);

BUFG bufg_adc_clk    (.O (adc_clk   ), .I (pll_adc_clk   ));
BUFG bufg_dac_clk_1x (.O (dac_clk_1x), .I (pll_dac_clk_1x));
BUFG bufg_dac_clk_2x (.O (dac_clk_2x), .I (pll_dac_clk_2x));
BUFG bufg_dac_clk_2p (.O (dac_clk_2p), .I (pll_dac_clk_2p));
BUFG bufg_ser_clk    (.O (ser_clk   ), .I (pll_ser_clk   ));
BUFG bufg_pwm_clk    (.O (pwm_clk   ), .I (pll_pwm_clk   ));
*/


// ADC reset (active low) 
always @(posedge clk_adc_125mhz_000deg)
adc_rstn <=  frstn[0] &  pll_locked;

// DAC reset (active high)
always @(posedge clk_adc_125mhz_000deg)
dac_rst  <= ~frstn[0] | ~pll_locked;

// PWM reset (active low)
always @(posedge clk_adc_250mhz_000deg)
pwm_rstn <=  frstn[0] &  pll_locked;

////////////////////////////////////////////////////////////////////////////////
// ADC IO
////////////////////////////////////////////////////////////////////////////////

// generating ADC clock is disabled
assign adc_clk_o = 2'b10;
//ODDR i_adc_clk_p ( .Q(adc_clk_o[0]), .D1(1'b1), .D2(1'b0), .C(fclk[0]), .CE(1'b1), .R(1'b0), .S(1'b0));
//ODDR i_adc_clk_n ( .Q(adc_clk_o[1]), .D1(1'b0), .D2(1'b1), .C(fclk[0]), .CE(1'b1), .R(1'b0), .S(1'b0));

// ADC clock duty cycle stabilizer is enabled
assign adc_cdcs_o = 1'b1 ;

// IO block registers should be used here
// lowest 2 bits reserved for 16bit ADC
always @(posedge clk_adc_125mhz_000deg)
begin
  adc_dat_a <= adc_dat_a_i[16-1:2];
  adc_dat_b <= adc_dat_b_i[16-1:2];
end
    
// transform into 2's complement (negative slope)
assign adc_a = digital_loop ? dac_a : {adc_dat_a[14-1], ~adc_dat_a[14-2:0]};
assign adc_b = digital_loop ? dac_b : {adc_dat_b[14-1], ~adc_dat_b[14-2:0]};

////////////////////////////////////////////////////////////////////////////////
// DAC IO
////////////////////////////////////////////////////////////////////////////////

// Summation of ASG and PID signal perform saturation before sending to DAC 
assign dac_a_sum = asg_a + pid_a;
assign dac_b_sum = asg_b + pid_b;

// saturation
assign dac_a = (^dac_a_sum[15-1:15-2]) ? {dac_a_sum[15-1], {13{~dac_a_sum[15-1]}}} : dac_a_sum[14-1:0];
assign dac_b = (^dac_b_sum[15-1:15-2]) ? {dac_b_sum[15-1], {13{~dac_b_sum[15-1]}}} : dac_b_sum[14-1:0];

// output registers + signed to unsigned (also to negative slope)
always @(posedge clk_adc_125mhz_000deg)
begin
  dac_dat_a <= {dac_a[14-1], ~dac_a[14-2:0]};
  dac_dat_b <= {dac_b[14-1], ~dac_b[14-2:0]};
end

// DDR outputs
ODDR oddr_dac_clk          (.Q(dac_clk_o), .D1(1'b0     ), .D2(1'b1     ), .C(clk_adc_250mhz_315deg), .CE(1'b1), .R(dac_rst), .S(1'b0));
ODDR oddr_dac_wrt          (.Q(dac_wrt_o), .D1(1'b0     ), .D2(1'b1     ), .C(clk_adc_250mhz_000deg), .CE(1'b1), .R(dac_rst), .S(1'b0));
ODDR oddr_dac_sel          (.Q(dac_sel_o), .D1(1'b1     ), .D2(1'b0     ), .C(clk_adc_125mhz_000deg), .CE(1'b1), .R(dac_rst), .S(1'b0));
ODDR oddr_dac_rst          (.Q(dac_rst_o), .D1(dac_rst  ), .D2(dac_rst  ), .C(clk_adc_125mhz_000deg), .CE(1'b1), .R(1'b0   ), .S(1'b0));
ODDR oddr_dac_dat [14-1:0] (.Q(dac_dat_o), .D1(dac_dat_b), .D2(dac_dat_a), .C(clk_adc_125mhz_000deg), .CE(1'b1), .R(dac_rst), .S(1'b0));

//---------------------------------------------------------------------------------
//  House Keeping

wire  [  8-1: 0] exp_p_in , exp_n_in ;
wire  [  8-1: 0] exp_p_out, exp_n_out;
wire  [  8-1: 0] exp_p_dir, exp_n_dir;

red_pitaya_hk i_hk (
  // system signals
  .clk_i           (  clk_adc_125mhz_000deg      ),  // clock
  .rstn_i          (  adc_rstn                   ),  // reset - active low
  // LED
  .led_o           (  led_o                      ),  // LED output
  // global configuration
  .digital_loop    (  digital_loop               ),
  // Expansion connector
  .exp_p_dat_i     (  exp_p_in                   ),  // input data
  .exp_p_dat_o     (  exp_p_out                  ),  // output data
  .exp_p_dir_o     (  exp_p_dir                  ),  // 1-output enable
  .exp_n_dat_i     (  exp_n_in                   ),
  .exp_n_dat_o     (  exp_n_out                  ),
  .exp_n_dir_o     (  exp_n_dir                  ),
   // System bus
  .sys_addr        (  sys_addr                   ),  // address
  .sys_wdata       (  sys_wdata                  ),  // write data
  .sys_sel         (  sys_sel                    ),  // write byte select
  .sys_wen         (  sys_wen[0]                 ),  // write enable
  .sys_ren         (  sys_ren[0]                 ),  // read enable
  .sys_rdata       (  sys_rdata[ 0*32+:32]       ),  // read data
  .sys_err         (  sys_err[0]                 ),  // error indicator
  .sys_ack         (  sys_ack[0]                 )   // acknowledge signal
);

IOBUF i_iobufp [8-1:0] (.O(exp_p_in), .IO(exp_p_io), .I(exp_p_out), .T(~exp_p_dir) );
IOBUF i_iobufn [8-1:0] (.O(exp_n_in), .IO(exp_n_io), .I(exp_n_out), .T(~exp_n_dir) );

//---------------------------------------------------------------------------------
//  Oscilloscope application

wire trig_asg_out ;

red_pitaya_scope i_scope (
  // ADC
  .adc_a_i         (  adc_a                      ),  // CH 1
  .adc_b_i         (  adc_b                      ),  // CH 2
  .adc_clk_i       (  clk_adc_125mhz_000deg      ),  // clock
  .adc_rstn_i      (  adc_rstn                   ),  // reset - active low
  .trig_ext_i      (  exp_p_in[0]                ),  // external trigger
  .trig_asg_i      (  trig_asg_out               ),  // ASG trigger
  // two AXI masters - concatenated
  .axi_clk_o       ( {axi_clk   [1], axi_clk   [0]} ),  // global clock
  .axi_rstn_o      ( {axi_rstn  [1], axi_rstn  [0]} ),  // global reset
  .axi_waddr_o     ( {axi_waddr [1], axi_waddr [0]} ),  // system write address
  .axi_wdata_o     ( {axi_wdata [1], axi_wdata [0]} ),  // system write data
  .axi_wsel_o      ( {axi_wsel  [1], axi_wsel  [0]} ),  // system write byte select
  .axi_wvalid_o    ( {axi_wvalid[1], axi_wvalid[0]} ),  // system write data valid
  .axi_wlen_o      ( {axi_wlen  [1], axi_wlen  [0]} ),  // system write burst length
  .axi_wfixed_o    ( {axi_wfixed[1], axi_wfixed[0]} ),  // system write burst type (fixed / incremental)
  .axi_werr_i      ( {axi_werr  [1], axi_werr  [0]} ),  // system write error
  .axi_wrdy_i      ( {axi_wrdy  [1], axi_wrdy  [0]} ),  // system write ready
  // System bus
  .sys_addr        (  sys_addr                   ),  // address
  .sys_wdata       (  sys_wdata                  ),  // write data
  .sys_sel         (  sys_sel                    ),  // write byte select
  .sys_wen         (  sys_wen[1]                 ),  // write enable
  .sys_ren         (  sys_ren[1]                 ),  // read enable
  .sys_rdata       (  sys_rdata[ 1*32+:32]       ),  // read data
  .sys_err         (  sys_err[1]                 ),  // error indicator
  .sys_ack         (  sys_ack[1]                 )   // acknowledge signal
);

//---------------------------------------------------------------------------------
//  DAC arbitrary signal generator

red_pitaya_asg i_asg (
   // DAC
  .dac_a_o         (  asg_a                      ),  // CH 1
  .dac_b_o         (  asg_b                      ),  // CH 2
  .dac_clk_i       (  clk_adc_125mhz_000deg      ),  // clock
  .dac_rstn_i      (  adc_rstn                   ),  // reset - active low
  .trig_a_i        (  exp_p_in[0]                ),
  .trig_b_i        (  exp_p_in[0]                ),
  .trig_out_o      (  trig_asg_out               ),
  // System bus
  .sys_addr        (  sys_addr                   ),  // address
  .sys_wdata       (  sys_wdata                  ),  // write data
  .sys_sel         (  sys_sel                    ),  // write byte select
  .sys_wen         (  sys_wen[2]                 ),  // write enable
  .sys_ren         (  sys_ren[2]                 ),  // read enable
  .sys_rdata       (  sys_rdata[ 2*32+:32]       ),  // read data
  .sys_err         (  sys_err[2]                 ),  // error indicator
  .sys_ack         (  sys_ack[2]                 )   // acknowledge signal
);

//---------------------------------------------------------------------------------
//  MIMO PID controller

red_pitaya_pid i_pid (
   // signals
  .clk_i           (  clk_adc_125mhz_000deg      ),  // clock
  .rstn_i          (  adc_rstn                   ),  // reset - active low
  .dat_a_i         (  adc_a                      ),  // in 1
  .dat_b_i         (  adc_b                      ),  // in 2
  .dat_a_o         (  pid_a                      ),  // out 1
  .dat_b_o         (  pid_b                      ),  // out 2
  // System bus
  .sys_addr        (  sys_addr                   ),  // address
  .sys_wdata       (  sys_wdata                  ),  // write data
  .sys_sel         (  sys_sel                    ),  // write byte select
  .sys_wen         (  sys_wen[3]                 ),  // write enable
  .sys_ren         (  sys_ren[3]                 ),  // read enable
  .sys_rdata       (  sys_rdata[ 3*32+:32]       ),  // read data
  .sys_err         (  sys_err[3]                 ),  // error indicator
  .sys_ack         (  sys_ack[3]                 )   // acknowledge signal
);

//---------------------------------------------------------------------------------
//  Analog mixed signals
//  XADC and slow PWM DAC control

wire  [ 24-1: 0] pwm_cfg_a;
wire  [ 24-1: 0] pwm_cfg_b;
wire  [ 24-1: 0] pwm_cfg_c;
wire  [ 24-1: 0] pwm_cfg_d;

red_pitaya_ams i_ams (
   // power test
  .clk_i           (  clk_adc_125mhz_000deg      ),  // clock
  .rstn_i          (  adc_rstn                   ),  // reset - active low
  // PWM configuration
  .dac_a_o         (  pwm_cfg_a                  ),
  .dac_b_o         (  pwm_cfg_b                  ),
  .dac_c_o         (  pwm_cfg_c                  ),
  .dac_d_o         (  pwm_cfg_d                  ),
   // System bus
  .sys_addr        (  sys_addr                   ),  // address
  .sys_wdata       (  sys_wdata                  ),  // write data
  .sys_sel         (  sys_sel                    ),  // write byte select
  .sys_wen         (  sys_wen[4]                 ),  // write enable
  .sys_ren         (  sys_ren[4]                 ),  // read enable
  .sys_rdata       (  sys_rdata[ 4*32+:32]       ),  // read data
  .sys_err         (  sys_err[4]                 ),  // error indicator
  .sys_ack         (  sys_ack[4]                 )   // acknowledge signal
);

red_pitaya_pwm i_pwm [4-1:0] (
  // system signals
  .clk   (clk_adc_250mhz_000deg),
  .rstn  (pwm_rstn),
  // configuration
  .cfg   ({pwm_cfg_d, pwm_cfg_c, pwm_cfg_b, pwm_cfg_a}),
  // PWM outputs
  .pwm_o (dac_pwm_o),
  .pwm_s ()
);

//---------------------------------------------------------------------------------
//  Daisy chain
//  simple communication module

wire daisy_rx_rdy ;
wire dly_clk = fclk[3];                              // 200MHz clock from PS - used for IDELAY (optionaly)

red_pitaya_daisy i_daisy (
   // SATA connector
  .daisy_p_o       (  daisy_p_o                  ),  // line 1 is clock capable
  .daisy_n_o       (  daisy_n_o                  ),
  .daisy_p_i       (  daisy_p_i                  ),  // line 1 is clock capable
  .daisy_n_i       (  daisy_n_i                  ),
   // Data
  .ser_clk_i       (  clk_adc_250mhz_000deg      ),  // high speed serial
  .dly_clk_i       (  dly_clk                    ),  // delay clock
   // TX
  .par_clk_i       (  clk_adc_125mhz_000deg      ),  // data paralel clock
  .par_rstn_i      (  adc_rstn                   ),  // reset - active low
  .par_rdy_o       (  daisy_rx_rdy               ),
  .par_dv_i        (  daisy_rx_rdy               ),
  .par_dat_i       (  16'h1234                   ),
   // RX
  .par_clk_o       (                             ),
  .par_rstn_o      (                             ),
  .par_dv_o        (                             ),
  .par_dat_o       (                             ),

  .debug_o         (/*led_o*/                    ),
   // System bus
  .sys_clk_i       (  sys_clk                    ),  // clock
  .sys_rstn_i      (  sys_rstn                   ),  // reset - active low
  .sys_addr_i      (  sys_addr                   ),  // address
  .sys_wdata_i     (  sys_wdata                  ),  // write data
  .sys_sel_i       (  sys_sel                    ),  // write byte select
  .sys_wen_i       (  sys_wen[5]                 ),  // write enable
  .sys_ren_i       (  sys_ren[5]                 ),  // read enable
  .sys_rdata_o     (  sys_rdata[ 5*32+:32]       ),  // read data
  .sys_err_o       (  sys_err[5]                 ),  // error indicator
  .sys_ack_o       (  sys_ack[5]                 )   // acknowledge signal
);

//---------------------------------------------------------------------------------
//  RadioBox module

red_pitaya_radiobox i_radiobox (
  // ADC
  .clk_adc_125mhz  (  clk_adc_125mhz_000deg      ),  // clock 125 MHz
  .clk_adc_20mhz   (  clk_adc_20mhz_000deg       ),  // clock  20 MHz
  .adc_rstn_i      (  adc_rstn                   ),  // reset - active low
/*
  .adc_a_i         (  adc_a                      ),  // CH 1
  .adc_b_i         (  adc_b                      ),  // CH 2
  .trig_ext_i      (  exp_p_in[0]                ),  // external trigger
  .trig_asg_i      (  trig_asg_out               ),  // ASG trigger
*/

/*
  // AXI1 master                         // AXI0 master
  .axi1_clk_o      (  axi_clk   [1]  ),  .axi0_clk_o      (  axi_clk   [0]  ),
  .axi1_rstn_o     (  axi_rstn  [1]  ),  .axi0_rstn_o     (  axi_rstn  [0]  ),
  .axi1_waddr_o    (  axi_waddr [1]  ),  .axi0_waddr_o    (  axi_waddr [0]  ),
  .axi1_wdata_o    (  axi_wdata [1]  ),  .axi0_wdata_o    (  axi_wdata [0]  ),
  .axi1_wsel_o     (  axi_wsel  [1]  ),  .axi0_wsel_o     (  axi_wsel  [0]  ),
  .axi1_wvalid_o   (  axi_wvalid[1]  ),  .axi0_wvalid_o   (  axi_wvalid[0]  ),
  .axi1_wlen_o     (  axi_wlen  [1]  ),  .axi0_wlen_o     (  axi_wlen  [0]  ),
  .axi1_wfixed_o   (  axi_wfixed[1]  ),  .axi0_wfixed_o   (  axi_wfixed[0]  ),
  .axi1_werr_i     (  axi_werr  [1]  ),  .axi0_werr_i     (  axi_werr  [0]  ),
  .axi1_wrdy_i     (  axi_wrdy  [1]  ),  .axi0_wrdy_i     (  axi_wrdy  [0]  ),
*/

  // System bus
  .sys_addr        (  sys_addr                   ),  // address
  .sys_wdata       (  sys_wdata                  ),  // write data
  .sys_sel         (  sys_sel                    ),  // write byte select
  .sys_wen         (  sys_wen[6]                 ),  // write enable
  .sys_ren         (  sys_ren[6]                 ),  // read enable
  .sys_rdata       (  sys_rdata[ 6*32+:32]       ),  // read data
  .sys_err         (  sys_err[6]                 ),  // error indicator
  .sys_ack         (  sys_ack[6]                 )   // acknowledge signal
);

endmodule
